module Kartsuba_reducer(
    output [162:0] d,
    input [324:0] a
);

    assign d[7:0]       = a[7:0]    ^a[170:163] ^a[324:317] ^a[286:279] ^a[253:246];                                                                            
    assign d[8]         = a[8]      ^a[171]     ^a[287]     ^a[254];                                                                                            
    assign d[16:9]      = a[16:9]   ^a[179:172] ^a[170:163] ^a[324:317] ^a[295:288] ^a[286:279] ^a[262:255] ^a[253:246];                                        
    assign d[45:17]     = a[45:17]  ^a[208:180] ^a[199:171] ^a[324:296] ^a[315:287] ^a[291:263] ^a[282:254];                                                    
    assign d[46]        = a[46]     ^a[209]     ^a[200]     ^a[316]     ^a[292]     ^a[283];                                                                    
    assign d[54:47]     = a[54:47]  ^a[217:210] ^a[208:201] ^a[170:163] ^a[324:317] ^a[324:317] ^a[286:279] ^a[300:293] ^a[291:284] ^a[253:246];                
    assign d[78:55]     = a[78:55]  ^a[241:218] ^a[232:209] ^a[194:171] ^a[310:287] ^a[324:301] ^a[315:292] ^a[277:254];                                        
    assign d[79]        = a[79]     ^a[242]     ^a[233]     ^a[195]     ^a[311]     ^a[316]     ^a[278];                                                        
    assign d[87:80]     = a[87:80]  ^a[250:243] ^a[241:234] ^a[203:196] ^a[170:163] ^a[324:317] ^a[319:312] ^a[286:279] ^a[324:317] ^a[286:279] ^a[253:246];    
    assign d[92:88]     = a[92:88]  ^a[255:251] ^a[246:242] ^a[208:204] ^a[175:171] ^a[324:320] ^a[291:287] ^a[291:287] ^a[258:254];                            
    assign d[125:93]    = a[125:93] ^a[288:256] ^a[279:246] ^a[241:209] ^a[208:176] ^a[324:292] ^a[324:292] ^a[291:259];                                       
    assign d[158:126]   = a[158:126]^a[321:289] ^a[312:280] ^a[274:242] ^a[241:209] ^a[324:292];                                                                
    assign d[161:159]   = a[161:159]^a[324:322] ^a[315:313] ^a[277:275] ^a[244:242];                                                                            
    assign d[162]       = a[162]    ^a[316]     ^a[278]     ^a[245];                                                                                            

endmodule